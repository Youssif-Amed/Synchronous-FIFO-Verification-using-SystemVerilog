package shared_pkg;
    int correct_count = 0;
    int error_count   = 0;
    bit test_finished;
endpackage